module wires ( input [3:0]x,y,
output [7:0]z);
assign z=x*y;
endmodule